* RLC

vin vin 0 1.8 PULSE 0 1.8 1m 1m 1m 20 40

.op
R1 vin 1 2
L1 1 out 1
C1 out 0 1

.tran 1m 16 0

.end
