* RLC

Vin vin 0 1.8

R1 vin out 10k
L1 out 0 5n
C1 out 0 1p

.op
.op

.end
