* RC

vin vin 0 1.8 PULSE 0 1.8 1n 1n 1n 100n 200n

.op
R1 vin out 10k
C1 out 0 1p

.tran 1n 500n 0

.end
