* staticDCStamp.sp

R1 1 0 0.1
G2 1 0 1 2 20
R3 1 2 0.2 
R4 2 0 0.5
I5 0 2 1.2
V6 3 2 1.3
E7 0 4 2 1 30
R8 3 4 0.4

.op

.end
