*Parser Test 

error1_here

vdd vdd 0 1.8

R1 vdd 1 5k
error2_here
C1 1 0 500f
L1 1 ab 2n
R2 ab c 2
Ila c 0 1m

.end
