* RC

vin vin 0 1.8 ac 1

R1 vin out 10k
C1 out 0 1p

.ac dec 1 1 1G

.end
